module top_tb;
  timeunit 1ps;
  timeprecision 1ps;

  //--------------------------------------------------------------------------------
  // Some basic parameters.
  //--------------------------------------------------------------------------------
  int clock_period_ps = 10;
  int timeout = 10000; // in cycles

  //--------------------------------------------------------------------------------
  // Clock generation
  //--------------------------------------------------------------------------------
  bit clk;
  initial clk = 1'b1;
  always #(clock_period_ps) clk = ~clk;

  //--------------------------------------------------------------------------------
  // Reset
  //--------------------------------------------------------------------------------
  bit rst;
  initial begin
    rst <= 1'b1;
    repeat (10) @(posedge clk);
    rst <= 1'b0;
  end


  //--------------------------------------------------------------------------------
  // Timeout setup
  //--------------------------------------------------------------------------------
  always @(posedge clk) begin
    if (timeout == 0) begin
      $error("TB Error: Timed out");
      $finish;
    end
    timeout <= timeout - 1;
  end

  //--------------------------------------------------------------------------------
  // Wave dumping
  //--------------------------------------------------------------------------------
  initial begin
    $fsdbDumpfile("dump.fsdb");
    $fsdbDumpvars(0, "+all");
  end

  //--------------------------------------------------------------------------------
  // Signals to connect to DUT.
  //--------------------------------------------------------------------------------

  // TODO for you: put here the I/O signals for the DUT.

  //--------------------------------------------------------------------------------
  // DUT instance
  //--------------------------------------------------------------------------------

  // TODO for you: instantiate the DUT.


  //--------------------------------------------------------------------------------
  // Tasks for verification
  //--------------------------------------------------------------------------------

  // TODO for you: verify the tasks!

  // Hint:
  /* task verify_task0();
    @(posedge clk);
    assert (task0_q === '0) else ...;
    task0_d <= $urandom();
    // assert something about task0_q
  endtask : verify_task0 */


  //--------------------------------------------------------------------------------
  // Helper functions
  //--------------------------------------------------------------------------------
  function print_seperator();
    repeat (80) $write("=");
    $write("\n");
  endfunction : print_seperator


  //--------------------------------------------------------------------------------
  // Main process
  //--------------------------------------------------------------------------------
  initial begin
    print_seperator();
    $finish;
  end

  final begin
    print_seperator();
  end

endmodule
